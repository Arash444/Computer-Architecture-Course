module Or(input a,b,output w);
	assign w = a | b;
endmodule
