module TB();
	reg clkk=1,initt=1;
	MIPS UUT(clkk,initt);
	always#10 clkk = ~clkk;
	initial begin
		#20 initt = 0;
		#1000 $stop;
	end
endmodule