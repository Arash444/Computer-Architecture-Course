module And(input a,b,output w);
	assign w = a&b;
endmodule